--sumador completo adder4 usando funcion
package ldl_bib is

component decobin2hex7seg is
   port( 

    ent:in   bit_vector(3 downto 0);
    sal :out  bit_vector(6 downto 0)
	
       );
end component decobin2hex7seg ;

end package ldl_bib;


	
